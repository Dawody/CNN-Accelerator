LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;


PACKAGE PKG IS

SUBTYPE BYTE IS STD_LOGIC_VECTOR(7 DOWNTO 0);
SUBTYPE ADDRESS IS STD_LOGIC_VECTOR(16 DOWNTO 0);
type five_bytes is array (0 to 4) of BYTE;



END PKG;



